`default_nettype none
`timescale 1ns/1ns

module vga_demo(
    input clk,
    input reset,
    output vga_h_sync,
    output vga_v_sync,
    output reg[3:0] vga_r,
    output reg[3:0] vga_g,
    output reg[3:0] vga_b
);

    wire [9:0] h_readwire, v_readwire;
    wire drawing_pixels;
    wire [3:0] rcol;
    wire [3:0] gcol;
    wire [3:0] bcol;
    
    sphere_renderer spb(
        .clk(clk),
        .reset(reset),
        .compr_hrw(h_readwire[9:3]),
        .compr_vrw(v_readwire[9:3]),
        .colorv(rcol),
        .startv(1'b1),
        .starth(1'b1),
        .top(21'd1398100)
    );

    sphere_renderer spg(
        .clk(clk),
        .reset(reset),
        .compr_hrw(h_readwire[9:3]),
        .compr_vrw(v_readwire[9:3]),
        .colorv(gcol),
        .startv(1'b1),
        .starth(1'b0),
        .top(21'd838860)
    );

    sphere_renderer spr(
        .clk(clk),
        .reset(reset),
        .compr_hrw(h_readwire[9:3]),
        .compr_vrw(v_readwire[9:3]),
        .colorv(bcol),
        .startv(1'b0),
        .starth(1'b1),
        .top(21'd1048576)
    );

    wire [11:0] bstream;
    wire [11:0] background;
    wire [11:0] foreground;

    wire [11:0] final_stream;
    wire [5:0] sumr, sumg, sumb;
    wire fbit;
    wire fvalue;
    assign background = 12'b000000000000;
    assign sumr = fvalue ? 4'b1111 : rcol + background[3:0] > 15 ? 15 : rcol + background[3:0];
    assign sumg = fvalue ? 4'b1111 : gcol + background[7:4] > 15 ? 15 : gcol + background[7:4];
    assign sumb = fvalue ? 4'b1111 : bcol + background[11:8] > 15 ? 15 : bcol + background[11:8];
    
    assign fbit = (h_readwire > 10'd475) & (h_readwire < 10'd635) & (v_readwire > 10'd420) &  (v_readwire < 10'd480);
    wire [9:0] imtar;
    assign fvalue = (drawing_pixels & fbit) ? !imbus[v_readwire - 10'd410][10'd635 - h_readwire] : 1'b0;
    
    wire [161:0] imbus [80:0]; 

    assign imbus[0] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[1] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[2] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[3] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[4] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[5] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[6] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[7] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[8] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[9] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[10] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[11] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[12] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[13] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[14] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[15] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[16] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[17] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[18] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[19] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[20] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[21] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[22] = 160'b1111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[23] = 160'b1111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[24] = 160'b1111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[25] = 160'b1111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[26] = 160'b1111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[27] = 160'b1111111111111111000000000000000000000000000000111111111111111111111111111111111111111100000000000011100111111111110011111111111111111111111111111111111111111111;
    assign imbus[28] = 160'b1111111111111100000000000000000000000000000000001111111111111111111111110000000111111100000000000011100111111111110011111111111111111111111111111111111111111111;
    assign imbus[29] = 160'b1111111111111000000000000111111111110000000000000111111111111111111111000000000001111111111111000111100111111111111111111111111111111111111111111111111111111111;
    assign imbus[30] = 160'b1111111111111000000000011111111111111110000000000111111111111111111110000111100000111111111111001111100111111111111111111111111111111111111111111111111111111111;
    assign imbus[31] = 160'b1111111111110000000001111111111111111111100000000011111111111111111100011111111100011111111110011111100100000111110011111000001001111100000011111000000111111111;
    assign imbus[32] = 160'b1111111111100000000011111111111111111111110000000001111111111111111000111111111110011111111100011111100000000011110011110000000001111000000001110000000011111111;
    assign imbus[33] = 160'b1111111111000000000000000000000001111111111000000000111111111111111001110000000110001111111000111111100001100011110011100001100001110000110000110001110011111111;
    assign imbus[34] = 160'b1111111111000000000000000000000001111110011100000000111111111111110001100000000111001111110001111111100111110001110011100011110001110001111000110011111111111111;
    assign imbus[35] = 160'b1111111110000000000000000000000011111110011110000000011111111111110011100011000111001111110011111111100111110001110011100111111001110011111100110000111111111111;
    assign imbus[36] = 160'b1111111110000000000000000000000011111100011111000000011111111111110011100111100111001111100111111111100111110001110011100111111001110011111100111000000111111111;
    assign imbus[37] = 160'b1111111110000000111111111100000111111100011111000000011111111111110011100111100110001111000111111111100111110001110011100111111001110011111100111111000011111111;
    assign imbus[38] = 160'b1111111100000001111111111100000111111000011111100000001111111111110011100011000000011110001111111111100111110001110011100011110001110001111000111111110001111111;
    assign imbus[39] = 160'b1111111100000001111111111100001111111000001111100000001111111111110011100000000000111100011111111111100001100011110011100001100001110000110000110011100001111111;
    assign imbus[40] = 160'b1111111100000011111111111000001111110000001111110000001111111111111001110000000001111100000000000011100000000011110011110000000001111000000001110000000011111111;
    assign imbus[41] = 160'b1111111000000011111111111000011111110000001111110000000111111111111000111111111111111100000000000011100100000111110011111000001001111100000011111000000111111111;
    assign imbus[42] = 160'b1111111000000011111111110000011111100000001111110000000111111111111100011111111001111111111111111111111111111111111111111111110001111111111111111111111111111111;
    assign imbus[43] = 160'b1111111000000111111111110000111111100000001111110000000111111111111110000111100001111111111111111111111111111111111111110011100001111111111111111111111111111111;
    assign imbus[44] = 160'b1111111000000111111111100000111111000000000111111000000111111111111111000000000011111111111111111111111111111111111111110000000011111111111111111111111111111111;
    assign imbus[45] = 160'b1111111000000111111111100001111111000010000111111000000111111111111111100000001111111111111111111111111111111111111111111000000111111111111111111111111111111111;
    assign imbus[46] = 160'b1111111000000111111111000001111110000010000111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[47] = 160'b1111111000000111111111000011111110000110000111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[48] = 160'b1111111000000111111110000011111100000111000011111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[49] = 160'b1111111000000011111110000111111100001111000011110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[50] = 160'b1111111000000011111100000111001000001111000011110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[51] = 160'b1111111100000011111100000000000000011111000011110000001111111111111000000011111111000001111110000000111111000000011111111111111111111111111111111111111111111111;
    assign imbus[52] = 160'b1111111100000011111000000000000000001111000011110000001111111111110000000001111110000000111100000000011110000000001111111111111111111111111111111111111111111111;
    assign imbus[53] = 160'b1111111100000001111000000000000000000001100001100000001111111111110001110000111100011000011100011100001110001110000111111111111111111111111111111111111111111111;
    assign imbus[54] = 160'b1111111100000001110000000000000000000111100001100000011111111111111111111000111100111100011111111110001111111111000111111111111111111111111111111111111111111111;
    assign imbus[55] = 160'b1111111110000000110000000000000001111111100001000000011111111111111111111000111000111110011111111110001111111111000111111111111111111111111111111111111111111111;
    assign imbus[56] = 160'b1111111110000000111111111000011011111111100000000000011111111111111111111000111000111110001111111110001111111111000111111111111111111111111111111111111111111111;
    assign imbus[57] = 160'b1111111111000000011111111111100011111111110000000000111111111111111111111001111000111110001111111110011111111111001111111111111111111111111111111111111111111111;
    assign imbus[58] = 160'b1111111111000000001111111110000011111111110000000000111111111111111111110011111000111110001111111100111111111110011111111111111111111111111111111111111111111111;
    assign imbus[59] = 160'b1111111111100000000111111110000111111111110000000001111111111111111111100011111000111110001111111000111111111100011111111111111111111111111111111111111111111111;
    assign imbus[60] = 160'b1111111111110000000011111100000111111111110000000011111111111111111111000111111000111110001111110001111111111000111111111111111111111111111111111111111111111111;
    assign imbus[61] = 160'b1111111111111000000000111100001111111111000000000111111111111111111110001111111000111110011111100011111111110001111111111111111111111111111111111111111111111111;
    assign imbus[62] = 160'b1111111111111100000000001000001111111100000000001111111111111111111100011111111100111100011111000111111111100011111111111111111111111111111111111111111111111111;
    assign imbus[63] = 160'b1111111111111110000000000000011111100000000000011111111111111111111000111111111100011000011110001111111111000111111111111111111111111111111111111111111111111111;
    assign imbus[64] = 160'b1111111111111111000000000000000000000000000000111111111111111111110000000000111110000000111100000000001110000000000111111111111111111111111111111111111111111111;
    assign imbus[65] = 160'b1111111111111111100000000000000000000000000001111111111111111111110000000000111111000001111100000000001110000000000111111111111111111111111111111111111111111111;
    assign imbus[66] = 160'b1111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[67] = 160'b1111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[68] = 160'b1111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[69] = 160'b1111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[70] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[71] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[72] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[73] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[74] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[75] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[76] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[77] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[78] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    assign imbus[79] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

    VGAcore core(
        .clk_25_175(clk),
        .reset(reset),
        .h_sync(vga_h_sync),
        .v_sync(vga_v_sync),
        .pixstream({sumr[3:0], sumg[3:0], sumb[3:0]}), //
        .hreadwire(h_readwire),
        .vreadwire(v_readwire),
        .drawing_pixels(drawing_pixels),
        .r(vga_r),
        .g(vga_g),
        .b(vga_b)
    );
endmodule
